 
* Copyright 2022 Mabrains
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT sky130_fd_pr__diode_pw2nd_05v5_lvt SUB
+ SUB D1_000_net_fail
+ SUB D1_001_net_fail
+ SUB D1_002_net_fail
+ SUB D1_003_net_fail
+ SUB D1_004_net_fail
+ SUB D1_005_net_fail
+ SUB D1_006_net_fail
+ SUB D1_007_net_fail
+ SUB D1_008_net_fail
+ SUB D1_009_net_fail
+ SUB D1_010_net_fail
+ SUB D1_011_net_fail
+ SUB D1_012_net_fail
+ SUB D1_013_net_fail
+ SUB D1_014_net_fail
+ SUB D1_015_net_fail
+ SUB D1_016_net_fail
+ SUB D1_017_net_fail
+ SUB D1_018_net_fail
+ SUB D1_019_net_fail
+ SUB D1_020_net_fail
+ SUB D1_021_net_fail
+ SUB D1_022_net_fail
+ SUB D1_023_net_fail
+ SUB D1_024_net_fail
+ SUB D1_025_net_fail
+ SUB D1_026_net_fail
+ SUB D1_027_net_fail
+ SUB D1_028_net_fail
+ SUB D1_029_net_fail
+ SUB D1_030_net_fail
+ SUB D1_031_net_fail
+ SUB D1_032_net_fail
+ SUB D1_033_net_fail
+ SUB D1_034_net_fail
+ SUB D1_035_net_fail
+ SUB D1_036_net_fail
+ SUB D1_037_net_fail
+ SUB D1_038_net_fail
+ SUB D1_039_net_fail
+ SUB D1_040_net_fail
+ SUB D1_041_net_fail
+ SUB D1_042_net_fail
+ SUB D1_043_net_fail
+ SUB D1_044_net_fail
+ SUB D1_045_net_fail
+ SUB D1_046_net_fail
+ SUB D1_047_net_fail
+ SUB D1_048_net_fail
+ SUB D1_049_net_fail
+ SUB D1_050_net_fail
+ SUB D1_051_net_fail
+ SUB D1_052_net_fail
+ SUB D1_053_net_fail
+ SUB D1_054_net_fail
+ SUB D1_055_net_fail
+ SUB D1_056_net_fail
+ SUB D1_057_net_fail
+ SUB D1_058_net_fail
+ SUB D1_059_net_fail
+ SUB D1_060_net_fail
+ SUB D1_061_net_fail
+ SUB D1_062_net_fail
+ SUB D1_063_net_fail

D000_net_fail SUB D1_000_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=0.24998625p P=2.2220999999999997u

D001_net_fail SUB D1_001_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=0.4999725p P=3.33315u

D002_net_fail SUB D1_002_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=0.74995875p P=4.4441999999999995u

D003_net_fail SUB D1_003_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=0.999945p P=5.55525u

D004_net_fail SUB D1_004_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=1.24993125p P=6.6663u

D005_net_fail SUB D1_005_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=1.4999175p P=7.777349999999999u

D006_net_fail SUB D1_006_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=1.7499037499999999p P=8.888399999999999u

D007_net_fail SUB D1_007_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=1.99989p P=9.99945u

D008_net_fail SUB D1_008_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=0.4999725p P=3.33315u

D009_net_fail SUB D1_009_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=0.999945p P=4.4441999999999995u

D010_net_fail SUB D1_010_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=1.4999175p P=5.55525u

D011_net_fail SUB D1_011_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=1.99989p P=6.6663u

D012_net_fail SUB D1_012_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=2.4998625p P=7.777349999999999u

D013_net_fail SUB D1_013_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=2.999835p P=8.888399999999999u

D014_net_fail SUB D1_014_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=3.4998074999999997p P=9.99945u

D015_net_fail SUB D1_015_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=3.99978p P=11.1105u

D016_net_fail SUB D1_016_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=0.74995875p P=4.4441999999999995u

D017_net_fail SUB D1_017_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=1.4999175p P=5.55525u

D018_net_fail SUB D1_018_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=2.24987625p P=6.6663u

D019_net_fail SUB D1_019_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=2.999835p P=7.777349999999999u

D020_net_fail SUB D1_020_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=3.74979375p P=8.888399999999999u

D021_net_fail SUB D1_021_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=4.4997525p P=9.99945u

D022_net_fail SUB D1_022_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=5.24971125p P=11.1105u

D023_net_fail SUB D1_023_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=5.99967p P=12.22155u

D024_net_fail SUB D1_024_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=0.999945p P=5.55525u

D025_net_fail SUB D1_025_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=1.99989p P=6.6663u

D026_net_fail SUB D1_026_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=2.999835p P=7.777349999999999u

D027_net_fail SUB D1_027_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=3.99978p P=8.888399999999999u

D028_net_fail SUB D1_028_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=4.999725p P=9.99945u

D029_net_fail SUB D1_029_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=5.99967p P=11.1105u

D030_net_fail SUB D1_030_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=6.9996149999999995p P=12.22155u

D031_net_fail SUB D1_031_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=7.99956p P=13.3326u

D032_net_fail SUB D1_032_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=1.24993125p P=6.6663u

D033_net_fail SUB D1_033_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=2.4998625p P=7.777349999999999u

D034_net_fail SUB D1_034_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=3.74979375p P=8.888399999999999u

D035_net_fail SUB D1_035_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=4.999725p P=9.99945u

D036_net_fail SUB D1_036_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=6.249656249999999p P=11.1105u

D037_net_fail SUB D1_037_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=7.4995875p P=12.22155u

D038_net_fail SUB D1_038_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=8.74951875p P=13.3326u

D039_net_fail SUB D1_039_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=9.99945p P=14.443649999999998u

D040_net_fail SUB D1_040_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=1.4999175p P=7.777349999999999u

D041_net_fail SUB D1_041_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=2.999835p P=8.888399999999999u

D042_net_fail SUB D1_042_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=4.4997525p P=9.99945u

D043_net_fail SUB D1_043_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=5.99967p P=11.1105u

D044_net_fail SUB D1_044_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=7.4995875p P=12.22155u

D045_net_fail SUB D1_045_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=8.999505p P=13.3326u

D046_net_fail SUB D1_046_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=10.4994225p P=14.443649999999998u

D047_net_fail SUB D1_047_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=11.99934p P=15.554699999999999u

D048_net_fail SUB D1_048_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=1.7499037499999999p P=8.888399999999999u

D049_net_fail SUB D1_049_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=3.4998074999999997p P=9.99945u

D050_net_fail SUB D1_050_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=5.24971125p P=11.1105u

D051_net_fail SUB D1_051_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=6.9996149999999995p P=12.22155u

D052_net_fail SUB D1_052_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=8.74951875p P=13.3326u

D053_net_fail SUB D1_053_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=10.4994225p P=14.443649999999998u

D054_net_fail SUB D1_054_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=12.24932625p P=15.554699999999999u

D055_net_fail SUB D1_055_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=13.999229999999999p P=16.66575u

D056_net_fail SUB D1_056_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=1.99989p P=9.99945u

D057_net_fail SUB D1_057_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=3.99978p P=11.1105u

D058_net_fail SUB D1_058_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=5.99967p P=12.22155u

D059_net_fail SUB D1_059_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=7.99956p P=13.3326u

D060_net_fail SUB D1_060_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=9.99945p P=14.443649999999998u

D061_net_fail SUB D1_061_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=11.99934p P=15.554699999999999u

D062_net_fail SUB D1_062_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=13.999229999999999p P=16.66575u

D063_net_fail SUB D1_063_net_fail sky130_fd_pr__diode_pw2nd_05v5_lvt A=15.99912p P=17.776799999999998u

.ENDS
 
* Copyright 2022 Mabrains
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT sky130_fd_pr__diode_pd2nw_05v5_lvt 
+ D0_000_lyr_fail D1_000_lyr_fail
+ D0_001_lyr_fail D1_001_lyr_fail
+ D0_002_lyr_fail D1_002_lyr_fail
+ D0_003_lyr_fail D1_003_lyr_fail
+ D0_004_lyr_fail D1_004_lyr_fail
+ D0_005_lyr_fail D1_005_lyr_fail
+ D0_006_lyr_fail D1_006_lyr_fail
+ D0_007_lyr_fail D1_007_lyr_fail
+ D0_008_lyr_fail D1_008_lyr_fail
+ D0_009_lyr_fail D1_009_lyr_fail
+ D0_010_lyr_fail D1_010_lyr_fail
+ D0_011_lyr_fail D1_011_lyr_fail
+ D0_012_lyr_fail D1_012_lyr_fail
+ D0_013_lyr_fail D1_013_lyr_fail
+ D0_014_lyr_fail D1_014_lyr_fail
+ D0_015_lyr_fail D1_015_lyr_fail
+ D0_016_lyr_fail D1_016_lyr_fail
+ D0_017_lyr_fail D1_017_lyr_fail
+ D0_018_lyr_fail D1_018_lyr_fail
+ D0_019_lyr_fail D1_019_lyr_fail
+ D0_020_lyr_fail D1_020_lyr_fail
+ D0_021_lyr_fail D1_021_lyr_fail
+ D0_022_lyr_fail D1_022_lyr_fail
+ D0_023_lyr_fail D1_023_lyr_fail
+ D0_024_lyr_fail D1_024_lyr_fail
+ D0_025_lyr_fail D1_025_lyr_fail
+ D0_026_lyr_fail D1_026_lyr_fail
+ D0_027_lyr_fail D1_027_lyr_fail
+ D0_028_lyr_fail D1_028_lyr_fail
+ D0_029_lyr_fail D1_029_lyr_fail
+ D0_030_lyr_fail D1_030_lyr_fail
+ D0_031_lyr_fail D1_031_lyr_fail
+ D0_032_lyr_fail D1_032_lyr_fail
+ D0_033_lyr_fail D1_033_lyr_fail
+ D0_034_lyr_fail D1_034_lyr_fail
+ D0_035_lyr_fail D1_035_lyr_fail
+ D0_036_lyr_fail D1_036_lyr_fail
+ D0_037_lyr_fail D1_037_lyr_fail
+ D0_038_lyr_fail D1_038_lyr_fail
+ D0_039_lyr_fail D1_039_lyr_fail
+ D0_040_lyr_fail D1_040_lyr_fail
+ D0_041_lyr_fail D1_041_lyr_fail
+ D0_042_lyr_fail D1_042_lyr_fail
+ D0_043_lyr_fail D1_043_lyr_fail
+ D0_044_lyr_fail D1_044_lyr_fail
+ D0_045_lyr_fail D1_045_lyr_fail
+ D0_046_lyr_fail D1_046_lyr_fail
+ D0_047_lyr_fail D1_047_lyr_fail
+ D0_048_lyr_fail D1_048_lyr_fail
+ D0_049_lyr_fail D1_049_lyr_fail
+ D0_050_lyr_fail D1_050_lyr_fail
+ D0_051_lyr_fail D1_051_lyr_fail
+ D0_052_lyr_fail D1_052_lyr_fail
+ D0_053_lyr_fail D1_053_lyr_fail
+ D0_054_lyr_fail D1_054_lyr_fail
+ D0_055_lyr_fail D1_055_lyr_fail
+ D0_056_lyr_fail D1_056_lyr_fail
+ D0_057_lyr_fail D1_057_lyr_fail
+ D0_058_lyr_fail D1_058_lyr_fail
+ D0_059_lyr_fail D1_059_lyr_fail
+ D0_060_lyr_fail D1_060_lyr_fail
+ D0_061_lyr_fail D1_061_lyr_fail
+ D0_062_lyr_fail D1_062_lyr_fail
+ D0_063_lyr_fail D1_063_lyr_fail

D000_lyr_fail D0_000_lyr_fail D1_000_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=0.2025p P=1.8u

D001_lyr_fail D0_001_lyr_fail D1_001_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=0.405p P=2.7u

D002_lyr_fail D0_002_lyr_fail D1_002_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=0.6075p P=3.6u

D003_lyr_fail D0_003_lyr_fail D1_003_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=0.81p P=4.5u

D004_lyr_fail D0_004_lyr_fail D1_004_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=1.0125p P=5.4u

D005_lyr_fail D0_005_lyr_fail D1_005_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=1.215p P=6.3u

D006_lyr_fail D0_006_lyr_fail D1_006_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=1.4175p P=7.2u

D007_lyr_fail D0_007_lyr_fail D1_007_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=1.62p P=8.1u

D008_lyr_fail D0_008_lyr_fail D1_008_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=0.405p P=2.7u

D009_lyr_fail D0_009_lyr_fail D1_009_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=0.81p P=3.6u

D010_lyr_fail D0_010_lyr_fail D1_010_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=1.215p P=4.5u

D011_lyr_fail D0_011_lyr_fail D1_011_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=1.62p P=5.4u

D012_lyr_fail D0_012_lyr_fail D1_012_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=2.025p P=6.3u

D013_lyr_fail D0_013_lyr_fail D1_013_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=2.43p P=7.2u

D014_lyr_fail D0_014_lyr_fail D1_014_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=2.835p P=8.1u

D015_lyr_fail D0_015_lyr_fail D1_015_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=3.24p P=9.0u

D016_lyr_fail D0_016_lyr_fail D1_016_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=0.6075p P=3.6u

D017_lyr_fail D0_017_lyr_fail D1_017_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=1.215p P=4.5u

D018_lyr_fail D0_018_lyr_fail D1_018_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=1.8225p P=5.4u

D019_lyr_fail D0_019_lyr_fail D1_019_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=2.43p P=6.3u

D020_lyr_fail D0_020_lyr_fail D1_020_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=3.0375p P=7.2u

D021_lyr_fail D0_021_lyr_fail D1_021_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=3.645p P=8.1u

D022_lyr_fail D0_022_lyr_fail D1_022_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=4.2525p P=9.0u

D023_lyr_fail D0_023_lyr_fail D1_023_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=4.86p P=9.9u

D024_lyr_fail D0_024_lyr_fail D1_024_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=0.81p P=4.5u

D025_lyr_fail D0_025_lyr_fail D1_025_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=1.62p P=5.4u

D026_lyr_fail D0_026_lyr_fail D1_026_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=2.43p P=6.3u

D027_lyr_fail D0_027_lyr_fail D1_027_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=3.24p P=7.2u

D028_lyr_fail D0_028_lyr_fail D1_028_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=4.05p P=8.1u

D029_lyr_fail D0_029_lyr_fail D1_029_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=4.86p P=9.0u

D030_lyr_fail D0_030_lyr_fail D1_030_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=5.67p P=9.9u

D031_lyr_fail D0_031_lyr_fail D1_031_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=6.48p P=10.8u

D032_lyr_fail D0_032_lyr_fail D1_032_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=1.0125p P=5.4u

D033_lyr_fail D0_033_lyr_fail D1_033_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=2.025p P=6.3u

D034_lyr_fail D0_034_lyr_fail D1_034_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=3.0375p P=7.2u

D035_lyr_fail D0_035_lyr_fail D1_035_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=4.05p P=8.1u

D036_lyr_fail D0_036_lyr_fail D1_036_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=5.0625p P=9.0u

D037_lyr_fail D0_037_lyr_fail D1_037_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=6.075p P=9.9u

D038_lyr_fail D0_038_lyr_fail D1_038_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=7.0875p P=10.8u

D039_lyr_fail D0_039_lyr_fail D1_039_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=8.1p P=11.7u

D040_lyr_fail D0_040_lyr_fail D1_040_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=1.215p P=6.3u

D041_lyr_fail D0_041_lyr_fail D1_041_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=2.43p P=7.2u

D042_lyr_fail D0_042_lyr_fail D1_042_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=3.645p P=8.1u

D043_lyr_fail D0_043_lyr_fail D1_043_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=4.86p P=9.0u

D044_lyr_fail D0_044_lyr_fail D1_044_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=6.075p P=9.9u

D045_lyr_fail D0_045_lyr_fail D1_045_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=7.29p P=10.8u

D046_lyr_fail D0_046_lyr_fail D1_046_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=8.505p P=11.7u

D047_lyr_fail D0_047_lyr_fail D1_047_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=9.72p P=12.6u

D048_lyr_fail D0_048_lyr_fail D1_048_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=1.4175p P=7.2u

D049_lyr_fail D0_049_lyr_fail D1_049_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=2.835p P=8.1u

D050_lyr_fail D0_050_lyr_fail D1_050_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=4.2525p P=9.0u

D051_lyr_fail D0_051_lyr_fail D1_051_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=5.67p P=9.9u

D052_lyr_fail D0_052_lyr_fail D1_052_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=7.0875p P=10.8u

D053_lyr_fail D0_053_lyr_fail D1_053_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=8.505p P=11.7u

D054_lyr_fail D0_054_lyr_fail D1_054_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=9.9225p P=12.6u

D055_lyr_fail D0_055_lyr_fail D1_055_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=11.34p P=13.5u

D056_lyr_fail D0_056_lyr_fail D1_056_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=1.62p P=8.1u

D057_lyr_fail D0_057_lyr_fail D1_057_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=3.24p P=9.0u

D058_lyr_fail D0_058_lyr_fail D1_058_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=4.86p P=9.9u

D059_lyr_fail D0_059_lyr_fail D1_059_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=6.48p P=10.8u

D060_lyr_fail D0_060_lyr_fail D1_060_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=8.1p P=11.7u

D061_lyr_fail D0_061_lyr_fail D1_061_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=9.72p P=12.6u

D062_lyr_fail D0_062_lyr_fail D1_062_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=11.34p P=13.5u

D063_lyr_fail D0_063_lyr_fail D1_063_lyr_fail sky130_fd_pr__diode_pd2nw_05v5_lvt A=12.96p P=14.4u

.ENDS
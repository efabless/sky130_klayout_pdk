 
* Copyright 2022 Mabrains
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT sky130_fd_pr__model__cap_mim_m4 
+ C0_000_lyr_fail C1_000_lyr_fail
+ C0_001_lyr_fail C1_001_lyr_fail
+ C0_002_lyr_fail C1_002_lyr_fail
+ C0_003_lyr_fail C1_003_lyr_fail
+ C0_004_lyr_fail C1_004_lyr_fail
+ C0_005_lyr_fail C1_005_lyr_fail
+ C0_006_lyr_fail C1_006_lyr_fail
+ C0_007_lyr_fail C1_007_lyr_fail
+ C0_008_lyr_fail C1_008_lyr_fail
+ C0_009_lyr_fail C1_009_lyr_fail
+ C0_010_lyr_fail C1_010_lyr_fail
+ C0_011_lyr_fail C1_011_lyr_fail
+ C0_012_lyr_fail C1_012_lyr_fail
+ C0_013_lyr_fail C1_013_lyr_fail
+ C0_014_lyr_fail C1_014_lyr_fail
+ C0_015_lyr_fail C1_015_lyr_fail
+ C0_016_lyr_fail C1_016_lyr_fail
+ C0_017_lyr_fail C1_017_lyr_fail
+ C0_018_lyr_fail C1_018_lyr_fail
+ C0_019_lyr_fail C1_019_lyr_fail
+ C0_020_lyr_fail C1_020_lyr_fail
+ C0_021_lyr_fail C1_021_lyr_fail
+ C0_022_lyr_fail C1_022_lyr_fail
+ C0_023_lyr_fail C1_023_lyr_fail
+ C0_024_lyr_fail C1_024_lyr_fail
+ C0_025_lyr_fail C1_025_lyr_fail
+ C0_026_lyr_fail C1_026_lyr_fail
+ C0_027_lyr_fail C1_027_lyr_fail
+ C0_028_lyr_fail C1_028_lyr_fail
+ C0_029_lyr_fail C1_029_lyr_fail
+ C0_030_lyr_fail C1_030_lyr_fail
+ C0_031_lyr_fail C1_031_lyr_fail
+ C0_032_lyr_fail C1_032_lyr_fail
+ C0_033_lyr_fail C1_033_lyr_fail
+ C0_034_lyr_fail C1_034_lyr_fail
+ C0_035_lyr_fail C1_035_lyr_fail
+ C0_036_lyr_fail C1_036_lyr_fail
+ C0_037_lyr_fail C1_037_lyr_fail
+ C0_038_lyr_fail C1_038_lyr_fail
+ C0_039_lyr_fail C1_039_lyr_fail
+ C0_040_lyr_fail C1_040_lyr_fail
+ C0_041_lyr_fail C1_041_lyr_fail
+ C0_042_lyr_fail C1_042_lyr_fail
+ C0_043_lyr_fail C1_043_lyr_fail
+ C0_044_lyr_fail C1_044_lyr_fail
+ C0_045_lyr_fail C1_045_lyr_fail
+ C0_046_lyr_fail C1_046_lyr_fail
+ C0_047_lyr_fail C1_047_lyr_fail
+ C0_048_lyr_fail C1_048_lyr_fail
+ C0_049_lyr_fail C1_049_lyr_fail
+ C0_050_lyr_fail C1_050_lyr_fail
+ C0_051_lyr_fail C1_051_lyr_fail
+ C0_052_lyr_fail C1_052_lyr_fail
+ C0_053_lyr_fail C1_053_lyr_fail
+ C0_054_lyr_fail C1_054_lyr_fail
+ C0_055_lyr_fail C1_055_lyr_fail
+ C0_056_lyr_fail C1_056_lyr_fail
+ C0_057_lyr_fail C1_057_lyr_fail
+ C0_058_lyr_fail C1_058_lyr_fail
+ C0_059_lyr_fail C1_059_lyr_fail
+ C0_060_lyr_fail C1_060_lyr_fail
+ C0_061_lyr_fail C1_061_lyr_fail
+ C0_062_lyr_fail C1_062_lyr_fail
+ C0_063_lyr_fail C1_063_lyr_fail
+ C0_064_lyr_fail C1_064_lyr_fail
+ C0_065_lyr_fail C1_065_lyr_fail
+ C0_066_lyr_fail C1_066_lyr_fail
+ C0_067_lyr_fail C1_067_lyr_fail
+ C0_068_lyr_fail C1_068_lyr_fail
+ C0_069_lyr_fail C1_069_lyr_fail
+ C0_070_lyr_fail C1_070_lyr_fail
+ C0_071_lyr_fail C1_071_lyr_fail
+ C0_072_lyr_fail C1_072_lyr_fail
+ C0_073_lyr_fail C1_073_lyr_fail
+ C0_074_lyr_fail C1_074_lyr_fail
+ C0_075_lyr_fail C1_075_lyr_fail
+ C0_076_lyr_fail C1_076_lyr_fail
+ C0_077_lyr_fail C1_077_lyr_fail
+ C0_078_lyr_fail C1_078_lyr_fail
+ C0_079_lyr_fail C1_079_lyr_fail
+ C0_080_lyr_fail C1_080_lyr_fail

C000_lyr_fail C0_000_lyr_fail C1_000_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=4p P=8u

C001_lyr_fail C0_001_lyr_fail C1_001_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=24p P=28u

C002_lyr_fail C0_002_lyr_fail C1_002_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=44p P=48u

C003_lyr_fail C0_003_lyr_fail C1_003_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=64p P=68u

C004_lyr_fail C0_004_lyr_fail C1_004_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=84p P=88u

C005_lyr_fail C0_005_lyr_fail C1_005_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=104p P=108u

C006_lyr_fail C0_006_lyr_fail C1_006_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=124p P=128u

C007_lyr_fail C0_007_lyr_fail C1_007_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=144p P=148u

C008_lyr_fail C0_008_lyr_fail C1_008_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=164p P=168u

C009_lyr_fail C0_009_lyr_fail C1_009_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=24p P=28u

C010_lyr_fail C0_010_lyr_fail C1_010_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=144p P=48u

C011_lyr_fail C0_011_lyr_fail C1_011_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=264p P=68u

C012_lyr_fail C0_012_lyr_fail C1_012_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=384p P=88u

C013_lyr_fail C0_013_lyr_fail C1_013_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=504p P=108u

C014_lyr_fail C0_014_lyr_fail C1_014_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=624p P=128u

C015_lyr_fail C0_015_lyr_fail C1_015_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=744p P=148u

C016_lyr_fail C0_016_lyr_fail C1_016_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=864p P=168u

C017_lyr_fail C0_017_lyr_fail C1_017_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=984p P=188u

C018_lyr_fail C0_018_lyr_fail C1_018_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=44p P=48u

C019_lyr_fail C0_019_lyr_fail C1_019_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=264p P=68u

C020_lyr_fail C0_020_lyr_fail C1_020_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=484p P=88u

C021_lyr_fail C0_021_lyr_fail C1_021_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=704p P=108u

C022_lyr_fail C0_022_lyr_fail C1_022_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=924p P=128u

C023_lyr_fail C0_023_lyr_fail C1_023_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=1144p P=148u

C024_lyr_fail C0_024_lyr_fail C1_024_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=1364p P=168u

C025_lyr_fail C0_025_lyr_fail C1_025_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=1584p P=188u

C026_lyr_fail C0_026_lyr_fail C1_026_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=1804p P=208u

C027_lyr_fail C0_027_lyr_fail C1_027_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=64p P=68u

C028_lyr_fail C0_028_lyr_fail C1_028_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=384p P=88u

C029_lyr_fail C0_029_lyr_fail C1_029_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=704p P=108u

C030_lyr_fail C0_030_lyr_fail C1_030_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=1024p P=128u

C031_lyr_fail C0_031_lyr_fail C1_031_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=1344p P=148u

C032_lyr_fail C0_032_lyr_fail C1_032_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=1664p P=168u

C033_lyr_fail C0_033_lyr_fail C1_033_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=1984p P=188u

C034_lyr_fail C0_034_lyr_fail C1_034_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=2304p P=208u

C035_lyr_fail C0_035_lyr_fail C1_035_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=2624p P=228u

C036_lyr_fail C0_036_lyr_fail C1_036_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=84p P=88u

C037_lyr_fail C0_037_lyr_fail C1_037_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=504p P=108u

C038_lyr_fail C0_038_lyr_fail C1_038_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=924p P=128u

C039_lyr_fail C0_039_lyr_fail C1_039_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=1344p P=148u

C040_lyr_fail C0_040_lyr_fail C1_040_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=1764p P=168u

C041_lyr_fail C0_041_lyr_fail C1_041_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=2184p P=188u

C042_lyr_fail C0_042_lyr_fail C1_042_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=2604p P=208u

C043_lyr_fail C0_043_lyr_fail C1_043_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=3024p P=228u

C044_lyr_fail C0_044_lyr_fail C1_044_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=3444p P=248u

C045_lyr_fail C0_045_lyr_fail C1_045_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=104p P=108u

C046_lyr_fail C0_046_lyr_fail C1_046_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=624p P=128u

C047_lyr_fail C0_047_lyr_fail C1_047_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=1144p P=148u

C048_lyr_fail C0_048_lyr_fail C1_048_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=1664p P=168u

C049_lyr_fail C0_049_lyr_fail C1_049_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=2184p P=188u

C050_lyr_fail C0_050_lyr_fail C1_050_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=2704p P=208u

C051_lyr_fail C0_051_lyr_fail C1_051_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=3224p P=228u

C052_lyr_fail C0_052_lyr_fail C1_052_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=3744p P=248u

C053_lyr_fail C0_053_lyr_fail C1_053_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=4264p P=268u

C054_lyr_fail C0_054_lyr_fail C1_054_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=124p P=128u

C055_lyr_fail C0_055_lyr_fail C1_055_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=744p P=148u

C056_lyr_fail C0_056_lyr_fail C1_056_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=1364p P=168u

C057_lyr_fail C0_057_lyr_fail C1_057_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=1984p P=188u

C058_lyr_fail C0_058_lyr_fail C1_058_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=2604p P=208u

C059_lyr_fail C0_059_lyr_fail C1_059_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=3224p P=228u

C060_lyr_fail C0_060_lyr_fail C1_060_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=3844p P=248u

C061_lyr_fail C0_061_lyr_fail C1_061_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=4464p P=268u

C062_lyr_fail C0_062_lyr_fail C1_062_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=5084p P=288u

C063_lyr_fail C0_063_lyr_fail C1_063_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=144p P=148u

C064_lyr_fail C0_064_lyr_fail C1_064_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=864p P=168u

C065_lyr_fail C0_065_lyr_fail C1_065_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=1584p P=188u

C066_lyr_fail C0_066_lyr_fail C1_066_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=2304p P=208u

C067_lyr_fail C0_067_lyr_fail C1_067_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=3024p P=228u

C068_lyr_fail C0_068_lyr_fail C1_068_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=3744p P=248u

C069_lyr_fail C0_069_lyr_fail C1_069_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=4464p P=268u

C070_lyr_fail C0_070_lyr_fail C1_070_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=5184p P=288u

C071_lyr_fail C0_071_lyr_fail C1_071_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=5904p P=308u

C072_lyr_fail C0_072_lyr_fail C1_072_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=164p P=168u

C073_lyr_fail C0_073_lyr_fail C1_073_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=984p P=188u

C074_lyr_fail C0_074_lyr_fail C1_074_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=1804p P=208u

C075_lyr_fail C0_075_lyr_fail C1_075_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=2624p P=228u

C076_lyr_fail C0_076_lyr_fail C1_076_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=3444p P=248u

C077_lyr_fail C0_077_lyr_fail C1_077_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=4264p P=268u

C078_lyr_fail C0_078_lyr_fail C1_078_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=5084p P=288u

C079_lyr_fail C0_079_lyr_fail C1_079_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=5904p P=308u

C080_lyr_fail C0_080_lyr_fail C1_080_lyr_fail sky130_fd_pr__model__cap_mim_m4 A=6724p P=328u

.ENDS
 
* Copyright 2022 Mabrains
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT sky130_fd_pr__res_iso_pw SUBSTRATE
+ R0_000_lyr_fail R1_000_lyr_fail
+ R0_001_lyr_fail R1_001_lyr_fail
+ R0_002_lyr_fail R1_002_lyr_fail
+ R0_003_lyr_fail R1_003_lyr_fail
+ R0_004_lyr_fail R1_004_lyr_fail
+ R0_005_lyr_fail R1_005_lyr_fail
+ R0_006_lyr_fail R1_006_lyr_fail
+ R0_007_lyr_fail R1_007_lyr_fail
+ R0_008_lyr_fail R1_008_lyr_fail
+ R0_009_lyr_fail R1_009_lyr_fail
+ R0_010_lyr_fail R1_010_lyr_fail
+ R0_011_lyr_fail R1_011_lyr_fail
+ R0_012_lyr_fail R1_012_lyr_fail
+ R0_013_lyr_fail R1_013_lyr_fail
+ R0_014_lyr_fail R1_014_lyr_fail
+ R0_015_lyr_fail R1_015_lyr_fail
+ R0_016_lyr_fail R1_016_lyr_fail
+ R0_017_lyr_fail R1_017_lyr_fail
+ R0_018_lyr_fail R1_018_lyr_fail
+ R0_019_lyr_fail R1_019_lyr_fail
+ R0_020_lyr_fail R1_020_lyr_fail
+ R0_021_lyr_fail R1_021_lyr_fail
+ R0_022_lyr_fail R1_022_lyr_fail
+ R0_023_lyr_fail R1_023_lyr_fail
+ R0_024_lyr_fail R1_024_lyr_fail
+ R0_025_lyr_fail R1_025_lyr_fail
+ R0_026_lyr_fail R1_026_lyr_fail
+ R0_027_lyr_fail R1_027_lyr_fail
+ R0_028_lyr_fail R1_028_lyr_fail
+ R0_029_lyr_fail R1_029_lyr_fail
+ R0_030_lyr_fail R1_030_lyr_fail
+ R0_031_lyr_fail R1_031_lyr_fail
+ R0_032_lyr_fail R1_032_lyr_fail
+ R0_033_lyr_fail R1_033_lyr_fail
+ R0_034_lyr_fail R1_034_lyr_fail
+ R0_035_lyr_fail R1_035_lyr_fail
+ R0_036_lyr_fail R1_036_lyr_fail
+ R0_037_lyr_fail R1_037_lyr_fail
+ R0_038_lyr_fail R1_038_lyr_fail
+ R0_039_lyr_fail R1_039_lyr_fail
+ R0_040_lyr_fail R1_040_lyr_fail
+ R0_041_lyr_fail R1_041_lyr_fail
+ R0_042_lyr_fail R1_042_lyr_fail
+ R0_043_lyr_fail R1_043_lyr_fail
+ R0_044_lyr_fail R1_044_lyr_fail
+ R0_045_lyr_fail R1_045_lyr_fail
+ R0_046_lyr_fail R1_046_lyr_fail
+ R0_047_lyr_fail R1_047_lyr_fail
+ R0_048_lyr_fail R1_048_lyr_fail
+ R0_049_lyr_fail R1_049_lyr_fail
+ R0_050_lyr_fail R1_050_lyr_fail
+ R0_051_lyr_fail R1_051_lyr_fail
+ R0_052_lyr_fail R1_052_lyr_fail
+ R0_053_lyr_fail R1_053_lyr_fail
+ R0_054_lyr_fail R1_054_lyr_fail
+ R0_055_lyr_fail R1_055_lyr_fail
+ R0_056_lyr_fail R1_056_lyr_fail
+ R0_057_lyr_fail R1_057_lyr_fail
+ R0_058_lyr_fail R1_058_lyr_fail
+ R0_059_lyr_fail R1_059_lyr_fail
+ R0_060_lyr_fail R1_060_lyr_fail
+ R0_061_lyr_fail R1_061_lyr_fail
+ R0_062_lyr_fail R1_062_lyr_fail
+ R0_063_lyr_fail R1_063_lyr_fail

R000_lyr_fail R0_000_lyr_fail R1_000_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=26.5u w=2.65u

R001_lyr_fail R0_001_lyr_fail R1_001_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=26.5u w=5.3u

R002_lyr_fail R0_002_lyr_fail R1_002_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=26.5u w=7.95u

R003_lyr_fail R0_003_lyr_fail R1_003_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=26.5u w=10.6u

R004_lyr_fail R0_004_lyr_fail R1_004_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=26.5u w=13.25u

R005_lyr_fail R0_005_lyr_fail R1_005_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=26.5u w=15.9u

R006_lyr_fail R0_006_lyr_fail R1_006_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=26.5u w=18.55u

R007_lyr_fail R0_007_lyr_fail R1_007_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=26.5u w=21.2u

R008_lyr_fail R0_008_lyr_fail R1_008_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=53.0u w=2.65u

R009_lyr_fail R0_009_lyr_fail R1_009_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=53.0u w=5.3u

R010_lyr_fail R0_010_lyr_fail R1_010_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=53.0u w=7.95u

R011_lyr_fail R0_011_lyr_fail R1_011_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=53.0u w=10.6u

R012_lyr_fail R0_012_lyr_fail R1_012_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=53.0u w=13.25u

R013_lyr_fail R0_013_lyr_fail R1_013_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=53.0u w=15.9u

R014_lyr_fail R0_014_lyr_fail R1_014_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=53.0u w=18.55u

R015_lyr_fail R0_015_lyr_fail R1_015_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=53.0u w=21.2u

R016_lyr_fail R0_016_lyr_fail R1_016_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=79.5u w=2.65u

R017_lyr_fail R0_017_lyr_fail R1_017_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=79.5u w=5.3u

R018_lyr_fail R0_018_lyr_fail R1_018_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=79.5u w=7.95u

R019_lyr_fail R0_019_lyr_fail R1_019_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=79.5u w=10.6u

R020_lyr_fail R0_020_lyr_fail R1_020_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=79.5u w=13.25u

R021_lyr_fail R0_021_lyr_fail R1_021_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=79.5u w=15.9u

R022_lyr_fail R0_022_lyr_fail R1_022_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=79.5u w=18.55u

R023_lyr_fail R0_023_lyr_fail R1_023_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=79.5u w=21.2u

R024_lyr_fail R0_024_lyr_fail R1_024_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=106.0u w=2.65u

R025_lyr_fail R0_025_lyr_fail R1_025_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=106.0u w=5.3u

R026_lyr_fail R0_026_lyr_fail R1_026_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=106.0u w=7.95u

R027_lyr_fail R0_027_lyr_fail R1_027_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=106.0u w=10.6u

R028_lyr_fail R0_028_lyr_fail R1_028_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=106.0u w=13.25u

R029_lyr_fail R0_029_lyr_fail R1_029_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=106.0u w=15.9u

R030_lyr_fail R0_030_lyr_fail R1_030_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=106.0u w=18.55u

R031_lyr_fail R0_031_lyr_fail R1_031_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=106.0u w=21.2u

R032_lyr_fail R0_032_lyr_fail R1_032_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=132.5u w=2.65u

R033_lyr_fail R0_033_lyr_fail R1_033_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=132.5u w=5.3u

R034_lyr_fail R0_034_lyr_fail R1_034_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=132.5u w=7.95u

R035_lyr_fail R0_035_lyr_fail R1_035_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=132.5u w=10.6u

R036_lyr_fail R0_036_lyr_fail R1_036_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=132.5u w=13.25u

R037_lyr_fail R0_037_lyr_fail R1_037_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=132.5u w=15.9u

R038_lyr_fail R0_038_lyr_fail R1_038_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=132.5u w=18.55u

R039_lyr_fail R0_039_lyr_fail R1_039_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=132.5u w=21.2u

R040_lyr_fail R0_040_lyr_fail R1_040_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=159.0u w=2.65u

R041_lyr_fail R0_041_lyr_fail R1_041_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=159.0u w=5.3u

R042_lyr_fail R0_042_lyr_fail R1_042_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=159.0u w=7.95u

R043_lyr_fail R0_043_lyr_fail R1_043_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=159.0u w=10.6u

R044_lyr_fail R0_044_lyr_fail R1_044_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=159.0u w=13.25u

R045_lyr_fail R0_045_lyr_fail R1_045_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=159.0u w=15.9u

R046_lyr_fail R0_046_lyr_fail R1_046_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=159.0u w=18.55u

R047_lyr_fail R0_047_lyr_fail R1_047_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=159.0u w=21.2u

R048_lyr_fail R0_048_lyr_fail R1_048_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=185.5u w=2.65u

R049_lyr_fail R0_049_lyr_fail R1_049_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=185.5u w=5.3u

R050_lyr_fail R0_050_lyr_fail R1_050_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=185.5u w=7.95u

R051_lyr_fail R0_051_lyr_fail R1_051_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=185.5u w=10.6u

R052_lyr_fail R0_052_lyr_fail R1_052_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=185.5u w=13.25u

R053_lyr_fail R0_053_lyr_fail R1_053_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=185.5u w=15.9u

R054_lyr_fail R0_054_lyr_fail R1_054_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=185.5u w=18.55u

R055_lyr_fail R0_055_lyr_fail R1_055_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=185.5u w=21.2u

R056_lyr_fail R0_056_lyr_fail R1_056_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=212.0u w=2.65u

R057_lyr_fail R0_057_lyr_fail R1_057_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=212.0u w=5.3u

R058_lyr_fail R0_058_lyr_fail R1_058_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=212.0u w=7.95u

R059_lyr_fail R0_059_lyr_fail R1_059_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=212.0u w=10.6u

R060_lyr_fail R0_060_lyr_fail R1_060_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=212.0u w=13.25u

R061_lyr_fail R0_061_lyr_fail R1_061_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=212.0u w=15.9u

R062_lyr_fail R0_062_lyr_fail R1_062_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=212.0u w=18.55u

R063_lyr_fail R0_063_lyr_fail R1_063_lyr_fail SUBSTRATE sky130_fd_pr__res_iso_pw l=212.0u w=21.2u

.ENDS
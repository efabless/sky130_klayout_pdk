 
* Copyright 2022 Mabrains
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT sky130_fd_pr__rf_npn_05v5_W1p00L4p00 C B E SUBSTRATE

Qx_lyr_fail C_lyr_fail B_lyr_fail E_lyr_fail SUBSTRATE sky130_fd_pr__rf_npn_05v5_W1p00L4p00

.ENDS
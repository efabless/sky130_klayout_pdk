 
* Copyright 2022 Mabrains
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT sky130_fd_pr__res_generic_po 
+ R0_000_net_fail R1_000_net_fail
+ R0_001_net_fail R1_001_net_fail
+ R0_002_net_fail R1_002_net_fail
+ R0_003_net_fail R1_003_net_fail
+ R0_004_net_fail R1_004_net_fail
+ R0_005_net_fail R1_005_net_fail
+ R0_006_net_fail R1_006_net_fail
+ R0_007_net_fail R1_007_net_fail
+ R0_008_net_fail R1_008_net_fail
+ R0_009_net_fail R1_009_net_fail
+ R0_010_net_fail R1_010_net_fail
+ R0_011_net_fail R1_011_net_fail
+ R0_012_net_fail R1_012_net_fail
+ R0_013_net_fail R1_013_net_fail
+ R0_014_net_fail R1_014_net_fail
+ R0_015_net_fail R1_015_net_fail
+ R0_016_net_fail R1_016_net_fail
+ R0_017_net_fail R1_017_net_fail
+ R0_018_net_fail R1_018_net_fail
+ R0_019_net_fail R1_019_net_fail
+ R0_020_net_fail R1_020_net_fail
+ R0_021_net_fail R1_021_net_fail
+ R0_022_net_fail R1_022_net_fail
+ R0_023_net_fail R1_023_net_fail
+ R0_024_net_fail R1_024_net_fail
+ R0_025_net_fail R1_025_net_fail
+ R0_026_net_fail R1_026_net_fail
+ R0_027_net_fail R1_027_net_fail
+ R0_028_net_fail R1_028_net_fail
+ R0_029_net_fail R1_029_net_fail
+ R0_030_net_fail R1_030_net_fail
+ R0_031_net_fail R1_031_net_fail
+ R0_032_net_fail R1_032_net_fail
+ R0_033_net_fail R1_033_net_fail
+ R0_034_net_fail R1_034_net_fail
+ R0_035_net_fail R1_035_net_fail
+ R0_036_net_fail R1_036_net_fail
+ R0_037_net_fail R1_037_net_fail
+ R0_038_net_fail R1_038_net_fail
+ R0_039_net_fail R1_039_net_fail
+ R0_040_net_fail R1_040_net_fail
+ R0_041_net_fail R1_041_net_fail
+ R0_042_net_fail R1_042_net_fail
+ R0_043_net_fail R1_043_net_fail
+ R0_044_net_fail R1_044_net_fail
+ R0_045_net_fail R1_045_net_fail
+ R0_046_net_fail R1_046_net_fail
+ R0_047_net_fail R1_047_net_fail
+ R0_048_net_fail R1_048_net_fail
+ R0_049_net_fail R1_049_net_fail
+ R0_050_net_fail R1_050_net_fail
+ R0_051_net_fail R1_051_net_fail
+ R0_052_net_fail R1_052_net_fail
+ R0_053_net_fail R1_053_net_fail
+ R0_054_net_fail R1_054_net_fail
+ R0_055_net_fail R1_055_net_fail
+ R0_056_net_fail R1_056_net_fail
+ R0_057_net_fail R1_057_net_fail
+ R0_058_net_fail R1_058_net_fail
+ R0_059_net_fail R1_059_net_fail
+ R0_060_net_fail R1_060_net_fail
+ R0_061_net_fail R1_061_net_fail
+ R0_062_net_fail R1_062_net_fail
+ R0_063_net_fail R1_063_net_fail

R000_net_fail R0_000_net_fail R1_000_net_fail sky130_fd_pr__res_generic_po l=2.0369249999999997u w=0.407385u

R001_net_fail R0_001_net_fail R1_001_net_fail sky130_fd_pr__res_generic_po l=2.0369249999999997u w=0.81477u

R002_net_fail R0_002_net_fail R1_002_net_fail sky130_fd_pr__res_generic_po l=2.0369249999999997u w=1.2221549999999999u

R003_net_fail R0_003_net_fail R1_003_net_fail sky130_fd_pr__res_generic_po l=2.0369249999999997u w=1.62954u

R004_net_fail R0_004_net_fail R1_004_net_fail sky130_fd_pr__res_generic_po l=2.0369249999999997u w=2.0369249999999997u

R005_net_fail R0_005_net_fail R1_005_net_fail sky130_fd_pr__res_generic_po l=2.0369249999999997u w=2.4443099999999998u

R006_net_fail R0_006_net_fail R1_006_net_fail sky130_fd_pr__res_generic_po l=2.0369249999999997u w=2.851695u

R007_net_fail R0_007_net_fail R1_007_net_fail sky130_fd_pr__res_generic_po l=2.0369249999999997u w=3.25908u

R008_net_fail R0_008_net_fail R1_008_net_fail sky130_fd_pr__res_generic_po l=4.073849999999999u w=0.407385u

R009_net_fail R0_009_net_fail R1_009_net_fail sky130_fd_pr__res_generic_po l=4.073849999999999u w=0.81477u

R010_net_fail R0_010_net_fail R1_010_net_fail sky130_fd_pr__res_generic_po l=4.073849999999999u w=1.2221549999999999u

R011_net_fail R0_011_net_fail R1_011_net_fail sky130_fd_pr__res_generic_po l=4.073849999999999u w=1.62954u

R012_net_fail R0_012_net_fail R1_012_net_fail sky130_fd_pr__res_generic_po l=4.073849999999999u w=2.0369249999999997u

R013_net_fail R0_013_net_fail R1_013_net_fail sky130_fd_pr__res_generic_po l=4.073849999999999u w=2.4443099999999998u

R014_net_fail R0_014_net_fail R1_014_net_fail sky130_fd_pr__res_generic_po l=4.073849999999999u w=2.851695u

R015_net_fail R0_015_net_fail R1_015_net_fail sky130_fd_pr__res_generic_po l=4.073849999999999u w=3.25908u

R016_net_fail R0_016_net_fail R1_016_net_fail sky130_fd_pr__res_generic_po l=6.110775u w=0.407385u

R017_net_fail R0_017_net_fail R1_017_net_fail sky130_fd_pr__res_generic_po l=6.110775u w=0.81477u

R018_net_fail R0_018_net_fail R1_018_net_fail sky130_fd_pr__res_generic_po l=6.110775u w=1.2221549999999999u

R019_net_fail R0_019_net_fail R1_019_net_fail sky130_fd_pr__res_generic_po l=6.110775u w=1.62954u

R020_net_fail R0_020_net_fail R1_020_net_fail sky130_fd_pr__res_generic_po l=6.110775u w=2.0369249999999997u

R021_net_fail R0_021_net_fail R1_021_net_fail sky130_fd_pr__res_generic_po l=6.110775u w=2.4443099999999998u

R022_net_fail R0_022_net_fail R1_022_net_fail sky130_fd_pr__res_generic_po l=6.110775u w=2.851695u

R023_net_fail R0_023_net_fail R1_023_net_fail sky130_fd_pr__res_generic_po l=6.110775u w=3.25908u

R024_net_fail R0_024_net_fail R1_024_net_fail sky130_fd_pr__res_generic_po l=8.147699999999999u w=0.407385u

R025_net_fail R0_025_net_fail R1_025_net_fail sky130_fd_pr__res_generic_po l=8.147699999999999u w=0.81477u

R026_net_fail R0_026_net_fail R1_026_net_fail sky130_fd_pr__res_generic_po l=8.147699999999999u w=1.2221549999999999u

R027_net_fail R0_027_net_fail R1_027_net_fail sky130_fd_pr__res_generic_po l=8.147699999999999u w=1.62954u

R028_net_fail R0_028_net_fail R1_028_net_fail sky130_fd_pr__res_generic_po l=8.147699999999999u w=2.0369249999999997u

R029_net_fail R0_029_net_fail R1_029_net_fail sky130_fd_pr__res_generic_po l=8.147699999999999u w=2.4443099999999998u

R030_net_fail R0_030_net_fail R1_030_net_fail sky130_fd_pr__res_generic_po l=8.147699999999999u w=2.851695u

R031_net_fail R0_031_net_fail R1_031_net_fail sky130_fd_pr__res_generic_po l=8.147699999999999u w=3.25908u

R032_net_fail R0_032_net_fail R1_032_net_fail sky130_fd_pr__res_generic_po l=10.184624999999999u w=0.407385u

R033_net_fail R0_033_net_fail R1_033_net_fail sky130_fd_pr__res_generic_po l=10.184624999999999u w=0.81477u

R034_net_fail R0_034_net_fail R1_034_net_fail sky130_fd_pr__res_generic_po l=10.184624999999999u w=1.2221549999999999u

R035_net_fail R0_035_net_fail R1_035_net_fail sky130_fd_pr__res_generic_po l=10.184624999999999u w=1.62954u

R036_net_fail R0_036_net_fail R1_036_net_fail sky130_fd_pr__res_generic_po l=10.184624999999999u w=2.0369249999999997u

R037_net_fail R0_037_net_fail R1_037_net_fail sky130_fd_pr__res_generic_po l=10.184624999999999u w=2.4443099999999998u

R038_net_fail R0_038_net_fail R1_038_net_fail sky130_fd_pr__res_generic_po l=10.184624999999999u w=2.851695u

R039_net_fail R0_039_net_fail R1_039_net_fail sky130_fd_pr__res_generic_po l=10.184624999999999u w=3.25908u

R040_net_fail R0_040_net_fail R1_040_net_fail sky130_fd_pr__res_generic_po l=12.22155u w=0.407385u

R041_net_fail R0_041_net_fail R1_041_net_fail sky130_fd_pr__res_generic_po l=12.22155u w=0.81477u

R042_net_fail R0_042_net_fail R1_042_net_fail sky130_fd_pr__res_generic_po l=12.22155u w=1.2221549999999999u

R043_net_fail R0_043_net_fail R1_043_net_fail sky130_fd_pr__res_generic_po l=12.22155u w=1.62954u

R044_net_fail R0_044_net_fail R1_044_net_fail sky130_fd_pr__res_generic_po l=12.22155u w=2.0369249999999997u

R045_net_fail R0_045_net_fail R1_045_net_fail sky130_fd_pr__res_generic_po l=12.22155u w=2.4443099999999998u

R046_net_fail R0_046_net_fail R1_046_net_fail sky130_fd_pr__res_generic_po l=12.22155u w=2.851695u

R047_net_fail R0_047_net_fail R1_047_net_fail sky130_fd_pr__res_generic_po l=12.22155u w=3.25908u

R048_net_fail R0_048_net_fail R1_048_net_fail sky130_fd_pr__res_generic_po l=14.258475u w=0.407385u

R049_net_fail R0_049_net_fail R1_049_net_fail sky130_fd_pr__res_generic_po l=14.258475u w=0.81477u

R050_net_fail R0_050_net_fail R1_050_net_fail sky130_fd_pr__res_generic_po l=14.258475u w=1.2221549999999999u

R051_net_fail R0_051_net_fail R1_051_net_fail sky130_fd_pr__res_generic_po l=14.258475u w=1.62954u

R052_net_fail R0_052_net_fail R1_052_net_fail sky130_fd_pr__res_generic_po l=14.258475u w=2.0369249999999997u

R053_net_fail R0_053_net_fail R1_053_net_fail sky130_fd_pr__res_generic_po l=14.258475u w=2.4443099999999998u

R054_net_fail R0_054_net_fail R1_054_net_fail sky130_fd_pr__res_generic_po l=14.258475u w=2.851695u

R055_net_fail R0_055_net_fail R1_055_net_fail sky130_fd_pr__res_generic_po l=14.258475u w=3.25908u

R056_net_fail R0_056_net_fail R1_056_net_fail sky130_fd_pr__res_generic_po l=16.295399999999997u w=0.407385u

R057_net_fail R0_057_net_fail R1_057_net_fail sky130_fd_pr__res_generic_po l=16.295399999999997u w=0.81477u

R058_net_fail R0_058_net_fail R1_058_net_fail sky130_fd_pr__res_generic_po l=16.295399999999997u w=1.2221549999999999u

R059_net_fail R0_059_net_fail R1_059_net_fail sky130_fd_pr__res_generic_po l=16.295399999999997u w=1.62954u

R060_net_fail R0_060_net_fail R1_060_net_fail sky130_fd_pr__res_generic_po l=16.295399999999997u w=2.0369249999999997u

R061_net_fail R0_061_net_fail R1_061_net_fail sky130_fd_pr__res_generic_po l=16.295399999999997u w=2.4443099999999998u

R062_net_fail R0_062_net_fail R1_062_net_fail sky130_fd_pr__res_generic_po l=16.295399999999997u w=2.851695u

R063_net_fail R0_063_net_fail R1_063_net_fail sky130_fd_pr__res_generic_po l=16.295399999999997u w=3.25908u

.ENDS